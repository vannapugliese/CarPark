`timescale 1ns / 100ps


module GlobalTime (

input wire clk;

output reg T;

);




endmodule